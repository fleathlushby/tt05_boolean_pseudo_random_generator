`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.09.2022 19:49:34
// Design Name: 
// Module Name: GF_MULS_4_shared
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// ------------------
//////////////////////////////////////////////////////////////////////////////////

(*keep = "true" , keep_hierarchy = "yes" *)
module GF_MULS_4_shared(input[3:0] in1_1, input[3:0] in1_2, input[3:0] in1_3, input[3:0] in2_1, input[3:0] in2_2, input[3:0] in2_3, output[3:0] out_1, output[3:0] out_2, output[3:0] out_3);

assign out_1[3] = ((in1_2[3] ^ in1_3[3]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[2] ^ in2_3[2])) ^((in1_2[3] ^ in1_3[3]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[0] ^ in2_3[0])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[0] ^ in2_3[0]));
assign out_2[3] = ((in1_1[3] & in2_3[3]) ^ (in2_1[3] & in1_3[3]) ^ (in1_1[3] & in2_1[3])) ^ ((in1_1[1] & in2_3[3]) ^ (in2_1[3] & in1_3[1]) ^ (in1_1[1] & in2_1[3])) ^ ((in1_1[0] & in2_3[3]) ^ (in2_1[3] & in1_3[0]) ^ (in1_1[0] & in2_1[3])) ^ ((in1_1[2] & in2_3[2]) ^ (in2_1[2] & in1_3[2]) ^ (in1_1[2] & in2_1[2])) ^ ((in1_1[1] & in2_3[2]) ^ (in2_1[2] & in1_3[1]) ^ (in1_1[1] & in2_1[2])) ^((in1_1[3] & in2_3[1]) ^ (in2_1[1] & in1_3[3]) ^ (in1_1[3] & in2_1[1])) ^ ((in1_1[2] & in2_3[1]) ^ (in2_1[1] & in1_3[2]) ^ (in1_1[2] & in2_1[1])) ^ ((in1_1[1] & in2_3[1]) ^ (in2_1[1] & in1_3[1]) ^ (in1_1[1] & in2_1[1])) ^ ((in1_1[0] & in2_3[1]) ^ (in2_1[1] & in1_3[0]) ^ (in1_1[0] & in2_1[1])) ^ ((in1_1[3] & in2_3[0]) ^ (in2_1[0] & in1_3[3]) ^ (in1_1[3] & in2_1[0])) ^ ((in1_1[1] & in2_3[0]) ^ (in2_1[0] & in1_3[1]) ^ (in1_1[1] & in2_1[0]));
assign out_3[3] = ((in1_1[3] & in2_2[3]) ^ (in2_1[3] & in1_2[3])) ^ ((in1_1[1] & in2_2[3]) ^ (in2_1[3] & in1_2[1])) ^ ((in1_1[0] & in2_2[3]) ^ (in2_1[3] & in1_2[0])) ^ ((in1_1[2] & in2_2[2]) ^ (in2_1[2] & in1_2[2])) ^ ((in1_1[1] & in2_2[2]) ^ (in2_1[2] & in1_2[1])) ^((in1_1[3] & in2_2[1]) ^ (in2_1[1] & in1_2[3])) ^ ((in1_1[2] & in2_2[1]) ^ (in2_1[1] & in1_2[2])) ^ ((in1_1[1] & in2_2[1]) ^ (in2_1[1] & in1_2[1])) ^ ((in1_1[0] & in2_2[1]) ^ (in2_1[1] & in1_2[0])) ^ ((in1_1[3] & in2_2[0]) ^ (in2_1[0] & in1_2[3])) ^ ((in1_1[1] & in2_2[0]) ^ (in2_1[0] & in1_2[1]));



assign out_1[2] = ((in1_2[2] ^ in1_3[2]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[2] ^ in2_3[2])) ^((in1_2[3] ^ in1_3[3]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[0] ^ in2_3[0])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[0] ^ in2_3[0]));
assign out_2[2] = ((in1_1[2] & in2_3[3]) ^ (in2_1[3] & in1_3[2]) ^ (in1_1[2] & in2_1[3])) ^ ((in1_1[1] & in2_3[3]) ^ (in2_1[3] & in1_3[1]) ^ (in1_1[1] & in2_1[3])) ^ ((in1_1[3] & in2_3[2]) ^ (in2_1[2] & in1_3[3]) ^ (in1_1[3] & in2_1[2])) ^ ((in1_1[2] & in2_3[2]) ^ (in2_1[2] & in1_3[2]) ^ (in1_1[2] & in2_1[2])) ^ ((in1_1[0] & in2_3[2]) ^ (in2_1[2] & in1_3[0]) ^ (in1_1[0] & in2_1[2])) ^((in1_1[3] & in2_3[1]) ^ (in2_1[1] & in1_3[3]) ^ (in1_1[3] & in2_1[1])) ^ ((in1_1[1] & in2_3[1]) ^ (in2_1[1] & in1_3[1]) ^ (in1_1[1] & in2_1[1])) ^ ((in1_1[2] & in2_3[0]) ^ (in2_1[0] & in1_3[2]) ^ (in1_1[2] & in2_1[0])) ^ ((in1_1[0] & in2_3[0]) ^ (in2_1[0] & in1_3[0]) ^ (in1_1[0] & in2_1[0]));
assign out_3[2] = ((in1_1[2] & in2_2[3]) ^ (in2_1[3] & in1_2[2])) ^ ((in1_1[1] & in2_2[3]) ^ (in2_1[3] & in1_2[1])) ^ ((in1_1[3] & in2_2[2]) ^ (in2_1[2] & in1_2[3])) ^ ((in1_1[2] & in2_2[2]) ^ (in2_1[2] & in1_2[2])) ^ ((in1_1[0] & in2_2[2]) ^ (in2_1[2] & in1_2[0])) ^ ((in1_1[3] & in2_2[1]) ^ (in2_1[1] & in1_2[3])) ^ ((in1_1[1] & in2_2[1]) ^ (in2_1[1] & in1_2[1])) ^ ((in1_1[2] & in2_2[0]) ^ (in2_1[0] & in1_2[2])) ^ ((in1_1[0] & in2_2[0]) ^ (in2_1[0] & in1_2[0]));



assign out_1[1] = ((in1_2[3] ^ in1_3[3]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[2] ^ in2_3[2])) ^((in1_2[1] ^ in1_3[1]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[0] ^ in2_3[0])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[0] ^ in2_3[0]));
assign out_2[1] = ((in1_1[3] & in2_3[3]) ^ (in2_1[3] & in1_3[3]) ^ (in1_1[3] & in2_1[3])) ^ ((in1_1[2] & in2_3[3]) ^ (in2_1[3] & in1_3[2]) ^ (in1_1[2] & in2_1[3])) ^ ((in1_1[1] & in2_3[3]) ^ (in2_1[3] & in1_3[1]) ^ (in1_1[1] & in2_1[3])) ^ ((in1_1[0] & in2_3[3]) ^ (in2_1[3] & in1_3[0]) ^ (in1_1[0] & in2_1[3])) ^ ((in1_1[3] & in2_3[2]) ^ (in2_1[2] & in1_3[3]) ^ (in1_1[3] & in2_1[2])) ^ ((in1_1[1] & in2_3[2]) ^ (in2_1[2] & in1_3[1]) ^ (in1_1[1] & in2_1[2])) ^ ((in1_1[3] & in2_3[1]) ^ (in2_1[1] & in1_3[3]) ^ (in1_1[3] & in2_1[1])) ^ ((in1_1[2] & in2_3[1]) ^ (in2_1[1] & in1_3[2]) ^ (in1_1[2] & in2_1[1])) ^ ((in1_1[1] & in2_3[1]) ^ (in2_1[1] & in1_3[1]) ^ (in1_1[1] & in2_1[1])) ^ ((in1_1[3] & in2_3[0]) ^ (in2_1[0] & in1_3[3]) ^ (in1_1[3] & in2_1[0])) ^ ((in1_1[0] & in2_3[0]) ^ (in2_1[0] & in1_3[0]) ^ (in1_1[0] & in2_1[0]));
assign out_3[1] = ((in1_1[3] & in2_2[3]) ^ (in2_1[3] & in1_2[3])) ^ ((in1_1[2] & in2_2[3]) ^ (in2_1[3] & in1_2[2])) ^ ((in1_1[1] & in2_2[3]) ^ (in2_1[3] & in1_2[1])) ^ ((in1_1[0] & in2_2[3]) ^ (in2_1[3] & in1_2[0])) ^ ((in1_1[3] & in2_2[2]) ^ (in2_1[2] & in1_2[3])) ^((in1_1[1] & in2_2[2]) ^ (in2_1[2] & in1_2[1])) ^ ((in1_1[3] & in2_2[1]) ^ (in2_1[1] & in1_2[3])) ^ ((in1_1[2] & in2_2[1]) ^ (in2_1[1] & in1_2[2])) ^ ((in1_1[1] & in2_2[1]) ^ (in2_1[1] & in1_2[1])) ^ ((in1_1[3] & in2_2[0]) ^ (in2_1[0] & in1_2[3])) ^ ((in1_1[0] & in2_2[0]) ^ (in2_1[0] & in1_2[0]));



assign out_1[0] = ((in1_2[3] ^ in1_3[3]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[3] ^ in2_3[3])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[2] ^ in2_3[2])) ^ ((in1_2[3] ^ in1_3[3]) & (in2_2[1] ^ in2_3[1])) ^((in1_2[0] ^ in1_3[0]) & (in2_2[1] ^ in2_3[1])) ^ ((in1_2[2] ^ in1_3[2]) & (in2_2[0] ^ in2_3[0])) ^ ((in1_2[1] ^ in1_3[1]) & (in2_2[0] ^ in2_3[0])) ^ ((in1_2[0] ^ in1_3[0]) & (in2_2[0] ^ in2_3[0]));
assign out_2[0] = ((in1_1[3] & in2_3[3]) ^ (in2_1[3] & in1_3[3]) ^ (in1_1[3] & in2_1[3])) ^ ((in1_1[1] & in2_3[3]) ^ (in2_1[3] & in1_3[1]) ^ (in1_1[1] & in2_1[3])) ^ ((in1_1[2] & in2_3[2]) ^ (in2_1[2] & in1_3[2]) ^ (in1_1[2] & in2_1[2])) ^ ((in1_1[0] & in2_3[2]) ^ (in2_1[2] & in1_3[0]) ^ (in1_1[0] & in2_1[2])) ^ ((in1_1[3] & in2_3[1]) ^ (in2_1[1] & in1_3[3]) ^ (in1_1[3] & in2_1[1])) ^((in1_1[0] & in2_3[1]) ^ (in2_1[1] & in1_3[0]) ^ (in1_1[0] & in2_1[1])) ^ ((in1_1[2] & in2_3[0]) ^ (in2_1[0] & in1_3[2]) ^ (in1_1[2] & in2_1[0])) ^ ((in1_1[1] & in2_3[0]) ^ (in2_1[0] & in1_3[1]) ^ (in1_1[1] & in2_1[0])) ^ ((in1_1[0] & in2_3[0]) ^ (in2_1[0] & in1_3[0]) ^ (in1_1[0] & in2_1[0]));
assign out_3[0] = ((in1_1[3] & in2_2[3]) ^ (in2_1[3] & in1_2[3])) ^ ((in1_1[1] & in2_2[3]) ^ (in2_1[3] & in1_2[1])) ^ ((in1_1[2] & in2_2[2]) ^ (in2_1[2] & in1_2[2])) ^ ((in1_1[0] & in2_2[2]) ^ (in2_1[2] & in1_2[0])) ^ ((in1_1[3] & in2_2[1]) ^ (in2_1[1] & in1_2[3])) ^((in1_1[0] & in2_2[1]) ^ (in2_1[1] & in1_2[0])) ^ ((in1_1[2] & in2_2[0]) ^ (in2_1[0] & in1_2[2])) ^ ((in1_1[1] & in2_2[0]) ^ (in2_1[0] & in1_2[1])) ^ ((in1_1[0] & in2_2[0]) ^ (in2_1[0] & in1_2[0]));

endmodule
