`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.09.2022 13:55:27
// Design Name: 
// Module Name: GF_INV_4_shared
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

(*keep = "true" , keep_hierarchy = "yes" *)
module GF_INV_4_shared(input[3:0] in_1, input[3:0] in_2, input[3:0] in_3, input[3:0] in_4, output[3:0] out_1, output[3:0] out_2, output[3:0] out_3, output[3:0] out_4);

assign out_1[3] = in_2[1] ^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ ((in_2[2] ^ in_3[2] ^ in_4[2]) & (in_2[1] ^ in_3[1] ^ in_4[1]) & (in_2[0] ^ in_3[0] ^ in_4[0]))
^ ((in_2[2] ^ in_3[2] ^ in_4[2]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ in_2[0];
assign out_2[3] = in_3[1] ^ ((in_1[3] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1])) ^ (in_1[2] & (in_3[1] ^ in_4[1]) & (in_3[0] ^ in_4[0])) ^ (in_1[1] &(in_3[2] ^ in_4[2]) & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[2] ^ in_4[2]) & (in_3[1] ^ in_4[1]))
^ (in_1[2] & in_1[1] & (in_3[0] ^ in_4[0])) ^ (in_1[2] & in_1[0] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & in_1[0] & (in_3[2] ^ in_4[2])) ^ (in_1[2] & in_1[1] & in_1[0])
^ (in_1[2] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[2] ^ in_4[2])) ^ (in_1[2] & in_1[1]) ^ in_3[0];
assign out_3[3] = in_4[1] ^ ((in_1[3] & in_2[1]) ^ (in_1[1] & in_2[3])) ^ (in_1[2] & in_1[1] & in_2[0]) ^ (in_1[2] & in_2[1] & in_1[0]) ^ (in_2[2] & in_1[1] & in_1[2]) ^ (in_1[2] & in_2[1] & in_2[0]) ^ (in_2[2] & in_1[1] & in_2[0]) ^ (in_2[2] & in_2[1] & in_1[0]) ^ (in_1[2] & in_2[1] & in_4[0])
^ (in_2[2] & in_1[1] & in_4[0]) ^ (in_1[2] & in_4[1] & in_2[0]) ^ (in_2[2] & in_4[1] & in_1[0]) ^ (in_4[2] & in_1[1] & in_2[0]) ^ (in_4[2] & in_2[1] & in_1[0]) ^ (in_1[2] & in_2[1]) ^ (in_1[1] & in_2[2]) ^ in_4[0];
assign out_4[3] = in_1[1] ^ (in_1[2] & in_2[1] & in_3[0]) ^ (in_1[2] & in_3[1] & in_2[0]) ^ (in_2[2] & in_1[1] & in_3[0]) ^ (in_2[2] & in_3[1] & in_1[0]) ^ (in_3[2] & in_1[1] & in_2[0]) ^ (in_3[2] & in_2[1] & in_1[0]) ^ in_1[0];


assign out_1[2] = ((in_2[2] ^ in_3[2] ^ in_4[2]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ ((in_2[2] ^ in_3[2] ^ in_4[2]) & (in_2[0] ^ in_3[0] ^ in_4[0])) ^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1]) & (in_2[0] ^ in_3[0] ^ in_4[0]))
^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ in_2[0];
assign out_2[2] = (in_1[2] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[2] ^ in_4[2])) ^ (in_1[2] & in_1[1]) ^ (in_1[2] & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[2] ^ in_4[2])) ^ (in_1[2] & in_1[0]) ^ (in_1[3] & (in_3[1] ^ in_4[1]) & (in_3[0] ^ in_4[0])) ^ (in_1[1] & (in_3[3] ^ in_4[3]) & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[3] ^ in_4[3]) & (in_3[1] ^ in_4[1]))
^ (in_1[3] & in_1[1] & (in_3[0] ^ in_4[0])) ^ (in_1[3] & in_1[0] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & in_1[0] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1] & in_1[0])
^ (in_1[3] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1]) ^ in_3[0];
assign out_3[2] = (in_1[2] & in_2[1]) ^ (in_1[1] & in_2[2]) ^ (in_1[2] & in_2[0]) ^ (in_1[0] & in_2[2]) ^ (in_1[3] & in_1[1] & in_2[0]) ^ (in_1[3] & in_2[1] & in_1[0]) ^ (in_2[3] & in_1[1] & in_1[3]) ^ (in_1[3] & in_2[1] & in_2[0]) ^ (in_2[3] & in_1[1] & in_2[0]) ^ (in_2[3] & in_2[1] & in_1[0]) ^ (in_1[3] & in_2[1] & in_4[0])
^ (in_2[3] & in_1[1] & in_4[0]) ^ (in_1[3] & in_4[1] & in_2[0]) ^ (in_2[3] & in_4[1] & in_1[0]) ^ (in_4[3] & in_1[1] & in_2[0]) ^ (in_4[3] & in_2[1] & in_1[0]) ^ (in_1[3] & in_2[1]) ^ (in_1[1] & in_2[3]) ^ in_4[0];
assign out_4[2] = (in_1[3] & in_2[1] & in_3[0]) ^ (in_1[3] & in_3[1] & in_2[0]) ^ (in_2[3] & in_1[1] & in_3[0]) ^ (in_2[3] & in_3[1] & in_1[0]) ^ (in_3[3] & in_1[1] & in_2[0]) ^ (in_3[3] & in_2[1] & in_1[0]) ^ in_1[0];


assign out_1[1] = in_1[3] ^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[0] ^ in_3[0] ^ in_4[0]) & (in_2[2] ^ in_3[2] ^ in_4[2]))
^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[0] ^ in_3[0] ^ in_4[0])) ^ in_2[2];
assign out_2[1] = in_2[3] ^ (in_1[3] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1]) ^ (in_1[3] & (in_3[0] ^ in_4[0]) & (in_3[2] ^ in_4[2])) ^ (in_1[0] & (in_3[3] ^ in_4[3]) & (in_3[2] ^ in_4[2])) ^ (in_1[2] & (in_3[3] ^ in_4[3]) & (in_3[0] ^ in_4[0]))
^ (in_1[3] & in_1[0] & (in_3[2] ^ in_4[2])) ^ (in_1[3] & in_1[2] & (in_3[0] ^ in_4[0])) ^ (in_1[0] & in_1[2] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[0] & in_1[2])
^ (in_1[3] & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[0]) ^ in_3[2];
assign out_3[1] = in_3[3] ^ (in_1[3] & in_2[1]) ^ (in_1[1] & in_2[3]) ^ (in_1[3] & in_1[0] & in_2[2]) ^ (in_1[3] & in_2[0] & in_1[2]) ^ (in_2[3] & in_1[0] & in_1[3]) ^ (in_1[3] & in_2[0] & in_2[2]) ^ (in_2[3] & in_1[0] & in_2[2]) ^ (in_2[3] & in_2[0] & in_1[2]) ^ (in_1[3] & in_2[0] & in_4[2])
^ (in_2[3] & in_1[0] & in_4[2]) ^ (in_1[3] & in_4[0] & in_2[2]) ^ (in_2[3] & in_4[0] & in_1[2]) ^ (in_4[3] & in_1[0] & in_2[2]) ^ (in_4[3] & in_2[0] & in_1[2]) ^ (in_1[3] & in_2[0]) ^ (in_1[0] & in_2[3]) ^ in_4[2];
assign out_4[1] = in_4[3] ^ (in_1[3] & in_2[0] & in_3[2]) ^ (in_1[3] & in_3[0] & in_2[2]) ^ (in_2[3] & in_1[0] & in_3[2]) ^ (in_2[3] & in_3[0] & in_1[2]) ^ (in_3[3] & in_1[0] & in_2[2]) ^ (in_3[3] & in_2[0] & in_1[2]) ^ 0 ^ in_1[2];



assign out_1[0] = ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[0] ^ in_3[0] ^ in_4[0])) ^ ((in_2[2] ^ in_3[2] ^ in_4[2]) & (in_2[0] ^ in_3[0] ^ in_4[0])) ^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1]) & (in_2[2] ^ in_3[2] ^ in_4[2]))
^ ((in_2[3] ^ in_3[3] ^ in_4[3]) & (in_2[1] ^ in_3[1] ^ in_4[1])) ^ in_2[2];
assign out_2[0] = (in_1[3] & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[0]) ^ (in_1[2] & (in_3[0] ^ in_4[0])) ^ (in_1[0] & (in_3[2] ^ in_4[2])) ^ (in_1[2] & in_1[0]) ^ (in_1[3] & (in_3[1] ^ in_4[1]) & (in_3[2] ^ in_4[2])) ^ (in_1[1] & (in_3[3] ^ in_4[3]) & (in_3[2] ^ in_4[2])) ^ (in_1[2] & (in_3[3] ^ in_4[3]) & (in_3[1] ^ in_4[1]))
^ (in_1[3] & in_1[1] & (in_3[2] ^ in_4[2])) ^ (in_1[3] & in_1[2] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & in_1[2] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1] & in_1[2])
^ (in_1[3] & (in_3[1] ^ in_4[1])) ^ (in_1[1] & (in_3[3] ^ in_4[3])) ^ (in_1[3] & in_1[1]) ^ in_3[2];
assign out_3[0] = (in_1[3] & in_2[0]) ^ (in_1[0] & in_2[3]) ^ (in_1[2] & in_2[0]) ^ (in_1[0] & in_2[2]) ^ (in_1[3] & in_1[1] & in_2[2]) ^ (in_1[3] & in_2[1] & in_1[2]) ^ (in_2[3] & in_1[1] & in_1[3]) ^ (in_1[3] & in_2[1] & in_2[2]) ^ (in_2[3] & in_1[1] & in_2[2]) ^ (in_2[3] & in_2[1] & in_1[2]) ^ (in_1[3] & in_2[1] & in_4[2])
^ (in_2[3] & in_1[1] & in_4[2]) ^ (in_1[3] & in_4[1] & in_2[2]) ^ (in_2[3] & in_4[1] & in_1[2]) ^ (in_4[3] & in_1[1] & in_2[2]) ^ (in_4[3] & in_2[1] & in_1[2]) ^ (in_1[3] & in_2[1]) ^ (in_1[1] & in_2[3]) ^ in_4[2];
assign out_4[0] = (in_1[3] & in_2[1] & in_3[2]) ^ (in_1[3] & in_3[1] & in_2[2]) ^ (in_2[3] & in_1[1] & in_3[2]) ^ (in_2[3] & in_3[1] & in_1[2]) ^ (in_3[3] & in_1[1] & in_2[2]) ^ (in_3[3] & in_2[1] & in_1[2]) ^ 0 ^ in_1[2];

endmodule
